.subckt INV_X1 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=14n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=10n TFIN=24n  HFIN=15n
.ends INV_X1

.subckt D_X1 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=14n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=10n TFIN=24n  HFIN=15n
.ends D_X1

.subckt INV_X2 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=27n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=20n TFIN=24n  HFIN=15n
.ends INV_X2

.subckt D_X2 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=27n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=20n TFIN=24n  HFIN=15n
.ends D_X2

.subckt INV_X3 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=40n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=30n TFIN=24n  HFIN=15n
.ends INV_X3

.subckt D_X3 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=40n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=30n TFIN=24n  HFIN=15n
.ends D_X3

.subckt INV_X4 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=52n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=40n TFIN=24n  HFIN=15n
.ends INV_X4

.subckt D_X4 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=52n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=40n TFIN=24n  HFIN=15n
.ends D_X4

.subckt INV_X5 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=64n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=50n TFIN=24n  HFIN=15n
.ends INV_X5

.subckt D_X5 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=64n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=50n TFIN=24n  HFIN=15n
.ends D_X5

.subckt INV_X6 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=77n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=60n TFIN=24n  HFIN=15n
.ends INV_X6

.subckt D_X6 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=77n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=60n TFIN=24n  HFIN=15n
.ends D_X6

.subckt INV_X7 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=89n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=70n TFIN=24n  HFIN=15n
.ends INV_X7

.subckt D_X7 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=89n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=70n TFIN=24n  HFIN=15n
.ends D_X7

.subckt INV_X8 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=101n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=80n TFIN=24n  HFIN=15n
.ends INV_X8

.subckt D_X8 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=101n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=80n TFIN=24n  HFIN=15n
.ends D_X8

.subckt INV_X9 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=114n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=90n TFIN=24n  HFIN=15n
.ends INV_X9

.subckt D_X9 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=114n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=90n TFIN=24n  HFIN=15n
.ends D_X9

.subckt INV_X10 VDD VSS A ZN
xmp1 ZN A VDD VDD pmos1 L=126n TFIN=24n  HFIN=15n
xmn1 ZN A VSS VSS nmos1 L=100n TFIN=24n  HFIN=15n
.ends INV_X10

.subckt D_X10 VDD VSS A 
xmp1 A A VDD VDD pmos1 L=126n TFIN=24n  HFIN=15n
xmn1 A A VSS VSS nmos1 L=100n TFIN=24n  HFIN=15n
.ends D_X10
